module u_top_z-top_z( );



endmodule
